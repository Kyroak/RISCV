--
-- VHDL Architecture RISCV_lib.dc_reg.behav
--
-- Created:
--          by - flxpuchr.meyer (pc032)
--          at - 15:55:37 05/16/23
--
-- using Mentor Graphics HDL Designer(TM) 2022.3 Built on 14 Jul 2022 at 13:56:12
--
library RISCV_lib;
USE RISCV_lib.opcode_word.ALL;
ARCHITECTURE behav OF dc_reg IS
BEGIN
    process(clk, res_n) is begin
   
    if res_n='0' then
      alu_mode_ex <= idle;
      value_a_1 <= (others => '0');
      reg_B_ex_1 <= (others => '0');
      imm_ex <= (others => '0');
      target_reg_ex <= (others => '0');
      fwd_sela_ex <= "00";
      fwd_selb_ex <= "00";
      fwd_selsd_ex <= '0';
            
      
      
  
    else
      if clk'event and clk = '1' then 
        alu_mode_ex   <= alu_mode_dc;
        value_a_1       <= reg_A_dc; 
        reg_B_ex_1      <= reg_B_dc; 
        imm_ex <= imm_bta_dc; 
        target_reg_ex <=  target_reg_dc;
        imm_to_alu_ex <= imm_to_alu_dc; 
        mem_mode_ex <= mem_mode_dc; 
        fwd_sela_ex <= fwd_sela_dc;
        fwd_selb_ex <= fwd_selb_dc;
        fwd_selsd_ex <= fwd_selsd_dc;
        
      end if;
    end if;
  end process;
END ARCHITECTURE behav;




