--
-- VHDL Architecture RISCV_lib.memory_control_unit_proofer.bahv
--
-- Created:
--          by - flxpuchr.meyer (pc032)
--          at - 17:39:30 06/20/23
--
-- using Mentor Graphics HDL Designer(TM) 2022.3 Built on 14 Jul 2022 at 13:56:12
--
ARCHITECTURE bahv OF memory_control_unit_proofer IS
BEGIN
END ARCHITECTURE bahv;

